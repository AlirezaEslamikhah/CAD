library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.Numeric_STD.ALL;

package pack is 
	type array8 is array(0 to 9) of std_logic_vector(0 to 7);
end pack;
