library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

package arr_package is
    type arr is array (0 to 7) of std_logic_vector(0 to 2);
end package arr_package;
